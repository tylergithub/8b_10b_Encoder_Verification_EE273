class msg;
	reg [9:0] dataout;
	reg [7:0] datain;
	reg pushin,startin,pushout,startout;
	
endclass
