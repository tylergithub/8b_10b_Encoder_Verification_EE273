// This is the output message class from the DUT:

class momsg;
	logic reset, startout, pushout;
	logic [8:0] dataout;
endclass