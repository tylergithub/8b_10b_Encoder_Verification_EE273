class mimsg;
	reg [9:0] dataout;
	reg [8:0] datain;
	reg pushin,startin,pushout,startout;
	
endclass
