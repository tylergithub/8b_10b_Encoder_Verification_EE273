// This is the output message class from the DUT:
// This class has not yet plug into the system yet
// I use this class for frame scoreboards: and data_frame_out_scoreboard
class momsg;
	logic reset, startout, pushout;
	logic [9:0] dataout;
endclass