// This is the input message class to the DUT:
// This class has not yet plug into the system yet
// I use this class for frame scoreboards: data_frame_in_scoreboard
class mimsg;
	logic reset, startin, pushin;
	logic [8:0] datain;
endclass