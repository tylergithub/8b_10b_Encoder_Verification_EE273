// This is the input message class to the DUT:

class mimsg;
	logic reset, startin, pushin;
	logic [8:0] datain;
endclass